library verilog;
use verilog.vl_types.all;
entity stimulus_counter is
end stimulus_counter;
