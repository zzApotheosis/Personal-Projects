library verilog;
use verilog.vl_types.all;
entity stimulus_seven_seg is
end stimulus_seven_seg;
