/*
 * Title: Test Module
 * Just testing how the button keys work.
 *
 * Date: 14 April 2017
 * Author: Steven Jennings
 * Copyright (C) 2017 Steven Jennings
 */

module Test(out, in);
	output out;
	input in;
	
	assign out = in;
endmodule
